//The drawback of ‘Ripple carry adder‘ is that it has a carry propagation delay that introduces slow computation.
//Since adders are used in designs like multipliers and divisions, it causes slowness in their computation. 
//To tackle this issue, a carry look-ahead adder (CLA) can be used that reduces propagation delay with additional hardware complexity

// https://vlsiverify.com/verilog/verilog-codes/carry-look-ahead-adder/

//CLA has introduced some functions like ‘carry generate (G)’ and ‘carry propagate (P)’ to boost the speed.
//Carry Generate (G): This function denotes how the carry is generated for single-bit two inputs regardless of any input carry.

//As we have seen in the full adder, carry is generated using the equation as A.B.
//Hence, G = A·B (similar to how carry is generated by full adder)
//Carry Propagate (P): This function denotes when the carry is propagated to the next stage with an addition whenever there is an input carry.

module CarryLookAheadAdder(
  input [3:0]A, B, 
  input Cin,
  output [3:0] S,
  output Cout
);
  wire [3:0] Ci; // Carry intermediate for intermediate computation
  
  assign Ci[0] = Cin;
  assign Ci[1] = (A[0] & B[0]) | ((A[0]^B[0]) & Ci[0]);
  //assign Ci[2] = (A[1] & B[1]) | ((A[1]^B[1]) & Ci[1]); expands to
  assign Ci[2] = (A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])));
  //assign Ci[3] = (A[2] & B[2]) | ((A[2]^B[2]) & Ci[2]); expands to
  assign Ci[3] = (A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))));
  //assign Cout  = (A[3] & B[3]) | ((A[3]^B[3]) & Ci[3]); expands to
  assign Cout  = (A[3] & B[3]) | ((A[3]^B[3]) & ((A[2] & B[2]) | ((A[2]^B[2]) & ((A[1] & B[1]) | ((A[1]^B[1]) & ((A[0] & B[0]) | ((A[0]^B[0]) & Ci[0])))))));

  assign S = A^B^Ci;
endmodule
